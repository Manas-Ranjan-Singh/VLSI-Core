//-------4bit_carry_lookhead_adder---------
//------------------ Half Adder ------------------
    module half_adder(
	                  g,
					   p,
					   a,
					   b);
	
    output              g;
    output              p;
    input               a;
    input               b;
	
    xor x1 (p, b, a);
    and a1 (g, b, a);
    endmodule

//------------------ XOR Gate ------------------
    module xor_gate(
    input i_cin,
    input i_pin,
    output o_sout
);
    xor x2 (o_sout, i_cin, i_pin);
endmodule

//------------------ Carry Look-Ahead Logic ------------------
    module addition(
    input [3:0] i_g,
    input [3:0] i_p,
    input       i_c,
    output[4:0] o_cout);
    assign o_cout[0] = i_c;
    assign o_cout[1] = i_g[0] | (i_p[0] & i_c);
    assign o_cout[2] = i_g[1] | (i_p[1] & i_g[0]) | (i_p[1] & i_p[0] & i_c);
    assign o_cout[3] = i_g[2] | (i_p[2] & i_g[1]) | (i_p[2] & i_p[1] & i_g[0]) | (i_p[2] & i_p[1] & i_p[0] & i_c);
    assign o_cout[4] = i_g[3] | (i_p[3] & i_g[2]) | (i_p[3] & i_p[2] & i_g[1]) |
                       (i_p[3] & i_p[2] & i_p[1] & i_g[0]) | (i_p[3] & i_p[2] & i_p[1] & i_p[0] & i_c);
    endmodule

//------------------ Main Module ------------------
module cla_4bit_add(
    output [3:0] o_s,
    output       o_c,
    input  [3:0] i_a,
    input  [3:0] i_b,
    input        i_cin
);
    wire [3:0] i_g;
    wire [3:0] i_p;
    wire [4:0] o_cout;

    // Half Adders for generate and propagate
    half_adder h0 (.g(i_g[0]),
                   .p(i_p[0]), 
                   .a(i_a[0]),
                   .b(i_b[0]));
    half_adder h1 (.g(i_g[1]),
                   .p(i_p[1]),
                   .a(i_a[1]),
                   .b(i_b[1]));
    half_adder h2 (.g(i_g[2]), 
                   .p(i_p[2]), 
                   .a(i_a[2]),
                   .b(i_b[2]));
    half_adder h3 (.g(i_g[3]),
                   .p(i_p[3]), 
                   .a(i_a[3]), 
                   .b(i_b[3]));

    // Carry Look-Ahead logic
    addition a1 (
                 .i_g(i_g),
                 .i_p(i_p),
                 .i_c(i_cin),
                 .o_cout(o_cout));

    // XOR gates for final sum output
    xor_gate x0 (.i_cin(o_cout[0]), 
                 .i_pin(i_p[0]), 
                 .o_sout(o_s[0]));
    xor_gate x1 (.i_cin(o_cout[1]), 
                 .i_pin(i_p[1]),
                 .o_sout(o_s[1]));
    xor_gate x2 (.i_cin(o_cout[2]), 
                 .i_pin(i_p[2]),
                 .o_sout(o_s[2]));
    xor_gate x3 (.i_cin(o_cout[3]),
                 .i_pin(i_p[3]),
                 .o_sout(o_s[3]));

    assign o_c = o_cout[4];

    endmodule
